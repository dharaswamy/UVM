interface adder_if;
  
  logic aclk,arst;
  logic [3:0] a,b;
  logic [4:0] y;
  
endinterface:adder_if