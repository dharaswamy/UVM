// Eda link : https://edaplayground.com/x/viML

// ( swamy ) please copy the code but don't change/modify the code here.

//=============================================================================================================================
// TOPIC NAME: UVM BASE CLASSES SOURCE CODES .

// i.uvm_drive
// ii.uvm_subscribe.

//=============================================================================================================================