interface sub_if;
  
  logic sclk,srst;
  logic [3:0] m,n;
  logic [4:0] z;
  
endinterface:sub_if