// Eda link : htt ps://edaplayground.com/x/JYPt 

// ( swamy ) please copy the code but don't change/modify the code here.

//===================================================================================================================
//     Topic Name: what is the "quasi static " in uvm
//===================================================================================================================

`include "uvm_macros.svh"
import uvm_pkg::*;
`include "user_component.sv"
`include "user_test.sv"

module tb;
  
  
  initial begin
  run_test("user_test");
  end
  
endmodule:tb